module LEGz_V3 (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4389593845 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(wire_16[7:0]), .en(wire_74), .out(arch_output_value));
  TC_Switch # (.UUID(64'd438959385 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_1 (.en(wire_29), .in(arch_input_value), .out(wire_51));
  TC_Program # (.UUID(64'd3388013681231061191 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_2F04A47E1BF0E0C7.w8.bin"), .ARG_SIG("Program_2F04A47E1BF0E0C7=%s")) Program_2 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_43 }), .out0(wire_101), .out1(wire_45), .out2(wire_42), .out3(wire_82));
  TC_Add # (.UUID(64'd1041402036361255287 ^ UUID), .BIT_WIDTH(64'd8)) Add8_3 (.in0(wire_1), .in1(wire_8), .ci(wire_23), .out(wire_80), .co());
  TC_And # (.UUID(64'd3149850418402764737 ^ UUID), .BIT_WIDTH(64'd8)) And8_4 (.in0(wire_1), .in1(wire_6), .out(wire_3));
  TC_Or # (.UUID(64'd2822446533483909240 ^ UUID), .BIT_WIDTH(64'd8)) Or8_5 (.in0(wire_1), .in1(wire_6), .out(wire_98));
  TC_Not # (.UUID(64'd3241827358460440603 ^ UUID), .BIT_WIDTH(64'd8)) Not8_6 (.in(wire_1), .out(wire_84));
  TC_Xor # (.UUID(64'd4419581709707773543 ^ UUID), .BIT_WIDTH(64'd8)) Xor8_7 (.in0(wire_1), .in1(wire_6), .out(wire_5));
  TC_Shr # (.UUID(64'd2969407248868243949 ^ UUID), .BIT_WIDTH(64'd8)) Shr8_8 (.in(wire_1), .shift(wire_6), .out(wire_53));
  TC_Shl # (.UUID(64'd4580910911811152089 ^ UUID), .BIT_WIDTH(64'd8)) Shl8_9 (.in(wire_1), .shift(wire_6), .out(wire_36));
  TC_Equal # (.UUID(64'd3366100765512475748 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_10 (.in0(wire_1), .in1(wire_6), .out(wire_35));
  TC_LessU # (.UUID(64'd1553277935616325458 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_11 (.in0(wire_1), .in1(wire_6), .out(wire_64));
  TC_Splitter8 # (.UUID(64'd418244241507724978 ^ UUID)) Splitter8_12 (.in(wire_45[7:0]), .out0(wire_38), .out1(wire_105), .out2(wire_103), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd2738989076623685468 ^ UUID)) Decoder3_13 (.dis(wire_65), .sel0(wire_38), .sel1(wire_105), .sel2(wire_103), .out0(wire_54), .out1(wire_87), .out2(wire_73), .out3(wire_97), .out4(wire_91), .out5(wire_22), .out6(wire_55), .out7(wire_31));
  TC_Counter # (.UUID(64'd2815704135892614591 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_14 (.clk(clk), .rst(rst), .save(wire_47), .in(wire_107), .out(wire_43));
  TC_Switch # (.UUID(64'd4540183510207418635 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_55), .in(wire_43), .out(wire_7_6));
  TC_Switch # (.UUID(64'd1066082560844542957 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_31), .in(wire_51), .out(wire_7_7));
  TC_Switch # (.UUID(64'd3167252235519358751 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_69), .in(wire_51), .out(wire_26_0));
  TC_Switch # (.UUID(64'd4014885166211024344 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_33), .in(wire_43), .out(wire_26_1));
  TC_Splitter8 # (.UUID(64'd1239159251500082281 ^ UUID)) Splitter8_19 (.in(wire_42[7:0]), .out0(wire_81), .out1(wire_110), .out2(wire_57), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd4136915607023856865 ^ UUID)) Decoder3_20 (.dis(wire_61), .sel0(wire_81), .sel1(wire_110), .sel2(wire_57), .out0(wire_52), .out1(wire_83), .out2(wire_85), .out3(wire_71), .out4(wire_104), .out5(wire_72), .out6(wire_33), .out7(wire_69));
  TC_Decoder3 # (.UUID(64'd1368739002161310908 ^ UUID)) Decoder3_21 (.dis(wire_63), .sel0(wire_14), .sel1(wire_79), .sel2(wire_0), .out0(wire_106), .out1(wire_99), .out2(wire_92), .out3(wire_50), .out4(wire_100), .out5(wire_25), .out6(wire_77), .out7(wire_74));
  TC_Splitter8 # (.UUID(64'd617943033813612701 ^ UUID)) Splitter8_22 (.in(wire_70), .out0(wire_14), .out1(wire_79), .out2(wire_0), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Or # (.UUID(64'd1925351272301252007 ^ UUID), .BIT_WIDTH(64'd1)) Or_23 (.in0(wire_31), .in1(wire_69), .out(wire_29));
  TC_Splitter8 # (.UUID(64'd2147155845543724529 ^ UUID)) Splitter8_24 (.in(wire_101[7:0]), .out0(wire_66), .out1(wire_56), .out2(wire_10), .out3(wire_12), .out4(wire_49), .out5(wire_30), .out6(wire_17), .out7(wire_20));
  TC_Or3 # (.UUID(64'd757853392458353090 ^ UUID), .BIT_WIDTH(64'd1)) Or3_25 (.in0(wire_12), .in1(wire_49), .in2(wire_30), .out(wire_11));
  TC_Decoder3 # (.UUID(64'd2003468714850951027 ^ UUID)) Decoder3_26 (.dis(wire_11), .sel0(wire_66), .sel1(wire_56), .sel2(wire_10), .out0(wire_34), .out1(wire_23), .out2(wire_93), .out3(wire_89), .out4(wire_2), .out5(wire_75), .out6(wire_68), .out7(wire_60));
  TC_Switch # (.UUID(64'd2253222201081204560 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_27 (.en(wire_34), .in(wire_6), .out(wire_8_1));
  TC_Switch # (.UUID(64'd147925994525832624 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_28 (.en(wire_23), .in(wire_94), .out(wire_8_0));
  TC_Switch # (.UUID(64'd4601921911051959516 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_29 (.en(wire_93), .in(wire_3), .out(wire_16_7[7:0]));
  TC_Switch # (.UUID(64'd4171828774110592372 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_30 (.en(wire_89), .in(wire_98), .out(wire_16_6[7:0]));
  TC_Switch # (.UUID(64'd1818751031091610596 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_31 (.en(wire_2), .in(wire_84), .out(wire_16_5[7:0]));
  TC_Switch # (.UUID(64'd432388317737828159 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_32 (.en(wire_75), .in(wire_5), .out(wire_16_4[7:0]));
  TC_Switch # (.UUID(64'd422541836763510756 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_33 (.en(wire_68), .in(wire_53), .out(wire_16_2[7:0]));
  TC_Switch # (.UUID(64'd4382418280579940787 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_34 (.en(wire_60), .in(wire_36), .out(wire_16_0[7:0]));
  TC_Switch # (.UUID(64'd757954125054826366 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_35 (.en(wire_40), .in(wire_80), .out(wire_16_8[7:0]));
  TC_Or # (.UUID(64'd225472282621155203 ^ UUID), .BIT_WIDTH(64'd1)) Or_36 (.in0(wire_23), .in1(wire_34), .out(wire_40));
  TC_Mux # (.UUID(64'd3280125520563703154 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_37 (.sel(wire_20), .in0(wire_7), .in1(wire_45[7:0]), .out(wire_1));
  TC_Mux # (.UUID(64'd3648217315728292116 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_38 (.sel(wire_17), .in0(wire_26), .in1(wire_42[7:0]), .out(wire_6));
  TC_Not # (.UUID(64'd1579709013959366529 ^ UUID), .BIT_WIDTH(64'd1)) Not_39 (.in(wire_35), .out(wire_59));
  TC_Switch # (.UUID(64'd1769265135327276709 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_40 (.en(wire_37), .in(wire_35), .out(wire_27_2));
  TC_Switch # (.UUID(64'd2122641125041326972 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_41 (.en(wire_76), .in(wire_59), .out(wire_27_0));
  TC_Switch # (.UUID(64'd1601096853491394715 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_42 (.en(wire_90), .in(wire_64), .out(wire_27_1));
  TC_Switch # (.UUID(64'd1078905049743716681 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_43 (.en(wire_102), .in(wire_96), .out(wire_27_3));
  TC_Switch # (.UUID(64'd1860793972291087573 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_44 (.en(wire_32), .in(wire_48), .out(wire_27_4));
  TC_Switch # (.UUID(64'd192072952801963368 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_45 (.en(wire_95), .in(wire_78), .out(wire_27_5));
  TC_Or # (.UUID(64'd1280724427812746177 ^ UUID), .BIT_WIDTH(64'd1)) Or_46 (.in0(wire_35), .in1(wire_64), .out(wire_96));
  TC_Not # (.UUID(64'd1812011019841672414 ^ UUID), .BIT_WIDTH(64'd1)) Not_47 (.in(wire_64), .out(wire_78));
  TC_And # (.UUID(64'd2746875659703072521 ^ UUID), .BIT_WIDTH(64'd1)) And_48 (.in0(wire_59), .in1(wire_78), .out(wire_48));
  TC_Decoder3 # (.UUID(64'd4406038464453274193 ^ UUID)) Decoder3_49 (.dis(wire_44), .sel0(wire_66), .sel1(wire_56), .sel2(wire_10), .out0(wire_37), .out1(wire_76), .out2(wire_90), .out3(wire_102), .out4(wire_32), .out5(wire_95), .out6(), .out7());
  TC_Not # (.UUID(64'd3752005200523597270 ^ UUID), .BIT_WIDTH(64'd1)) Not_50 (.in(wire_30), .out(wire_108));
  TC_Mux # (.UUID(64'd4485643867827663182 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_51 (.sel(wire_15), .in0(wire_16[7:0]), .in1(wire_88), .out(wire_107));
  TC_Or3 # (.UUID(64'd346060345491981688 ^ UUID), .BIT_WIDTH(64'd1)) Or3_52 (.in0(wire_108), .in1(wire_49), .in2(wire_12), .out(wire_44));
  TC_And # (.UUID(64'd2136258934406885543 ^ UUID), .BIT_WIDTH(64'd1)) And_53 (.in0(wire_4), .in1(wire_49), .out(wire_28));
  TC_And # (.UUID(64'd1672604342831427930 ^ UUID), .BIT_WIDTH(64'd1)) And_54 (.in0(wire_19), .in1(wire_49), .out(wire_39));
  TC_Decoder1 # (.UUID(64'd3203704870661654999 ^ UUID)) Decoder1_55 (.sel(wire_66), .out0(wire_4), .out1(wire_19));
  TC_Not # (.UUID(64'd4556354685172745997 ^ UUID), .BIT_WIDTH(64'd8)) Not8_56 (.in(wire_6), .out(wire_94));
  TC_Mux # (.UUID(64'd4437121133770719098 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_57 (.sel(wire_21), .in0(wire_82[7:0]), .in1(wire_45[7:0]), .out(wire_70));
  TC_Or # (.UUID(64'd3185911640361027442 ^ UUID), .BIT_WIDTH(64'd1)) Or_58 (.in0(wire_28), .in1(wire_46), .out(wire_21));
  TC_And # (.UUID(64'd1122576109677063165 ^ UUID), .BIT_WIDTH(64'd1)) And_59 (.in0(wire_12), .in1(wire_19), .out(wire_46));
  TC_And # (.UUID(64'd3520152224138576016 ^ UUID), .BIT_WIDTH(64'd1)) And_60 (.in0(wire_12), .in1(wire_4), .out(wire_67));
  TC_Or # (.UUID(64'd4325928675775570615 ^ UUID), .BIT_WIDTH(64'd1)) Or_61 (.in0(wire_67), .in1(wire_30), .out(wire_63));
  TC_Or # (.UUID(64'd4411131262145478365 ^ UUID), .BIT_WIDTH(64'd1)) Or_62 (.in0(wire_21), .in1(wire_20), .out(wire_65));
  TC_Or # (.UUID(64'd2446640561015928254 ^ UUID), .BIT_WIDTH(64'd1)) Or_63 (.in0(wire_21), .in1(wire_17), .out(wire_61));
  TC_Mux # (.UUID(64'd263177381119339096 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_64 (.sel(wire_41), .in0(wire_70), .in1(wire_45[7:0]), .out(wire_88));
  TC_Or3 # (.UUID(64'd1313293687935506487 ^ UUID), .BIT_WIDTH(64'd1)) Or3_65 (.in0(wire_15), .in1(wire_24), .in2(wire_77), .out(wire_47));
  TC_And # (.UUID(64'd4239975435082072874 ^ UUID), .BIT_WIDTH(64'd1)) And_66 (.in0(wire_30), .in1(wire_12), .out(wire_24));
  TC_And # (.UUID(64'd4171379149569873298 ^ UUID), .BIT_WIDTH(64'd1)) And_67 (.in0(wire_4), .in1(wire_24), .out(wire_41));
  TC_Add # (.UUID(64'd634203008895608581 ^ UUID), .BIT_WIDTH(64'd8)) Add8_68 (.in0(wire_43), .in1(wire_9), .ci(1'd0), .out(wire_62), .co());
  TC_Constant # (.UUID(64'd1557454806295191732 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_69 (.out(wire_9));
  TC_Mux # (.UUID(64'd2925228590958751190 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_70 (.sel(wire_41), .in0(wire_1), .in1(wire_62), .out(wire_58));
  TC_Or # (.UUID(64'd3489047166439471349 ^ UUID), .BIT_WIDTH(64'd1)) Or_71 (.in0(wire_67), .in1(wire_41), .out(wire_86));
  TC_Or # (.UUID(64'd3452358646011536940 ^ UUID), .BIT_WIDTH(64'd1)) Or_72 (.in0(wire_27), .in1(wire_41), .out(wire_15));
  TC_Or # (.UUID(64'd3985906689624227527 ^ UUID), .BIT_WIDTH(64'd1)) Or_73 (.in0(wire_109), .in1(wire_46), .out(wire_13));
  TC_And # (.UUID(64'd3665070101760230825 ^ UUID), .BIT_WIDTH(64'd1)) And_74 (.in0(wire_24), .in1(wire_19), .out(wire_109));
  TC_Ram # (.UUID(64'd657407049387028449 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_75 (.clk(clk), .rst(rst), .load(wire_28), .save(wire_39), .address({{24{1'b0}}, wire_18 }), .in0({{56{1'b0}}, wire_1 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_16_3), .out1(), .out2(), .out3());
  LegReg # (.UUID(64'd2211504464378337582 ^ UUID)) LegReg_76 (.clk(clk), .rst(rst), .Read_A(wire_54), .Read_B(wire_52), .Write(wire_106), .Write_Value(wire_16[7:0]), .Output_A(wire_7_0), .Output_B(wire_26_7), .Output());
  LegReg # (.UUID(64'd3273114815658507615 ^ UUID)) LegReg_77 (.clk(clk), .rst(rst), .Read_A(wire_22), .Read_B(wire_72), .Write(wire_25), .Write_Value(wire_16[7:0]), .Output_A(wire_7_5), .Output_B(wire_26_2), .Output(wire_18));
  STACK # (.UUID(64'd2648128136101199746 ^ UUID)) STACK_78 (.clk(clk), .rst(rst), .POP(wire_13), .PUSH(wire_86), .VALUE(wire_58), .OUTPUT(wire_16_1[7:0]));
  LegReg # (.UUID(64'd3220901936882606458 ^ UUID)) LegReg_79 (.clk(clk), .rst(rst), .Read_A(wire_91), .Read_B(wire_104), .Write(wire_100), .Write_Value(wire_16[7:0]), .Output_A(wire_7_4), .Output_B(wire_26_3), .Output());
  LegReg # (.UUID(64'd3301757283144249072 ^ UUID)) LegReg_80 (.clk(clk), .rst(rst), .Read_A(wire_97), .Read_B(wire_71), .Write(wire_50), .Write_Value(wire_16[7:0]), .Output_A(wire_7_3), .Output_B(wire_26_4), .Output());
  LegReg # (.UUID(64'd312975357935108921 ^ UUID)) LegReg_81 (.clk(clk), .rst(rst), .Read_A(wire_73), .Read_B(wire_85), .Write(wire_92), .Write_Value(wire_16[7:0]), .Output_A(wire_7_2), .Output_B(wire_26_5), .Output());
  LegReg # (.UUID(64'd3588865096648876778 ^ UUID)) LegReg_82 (.clk(clk), .rst(rst), .Read_A(wire_87), .Read_B(wire_83), .Write(wire_99), .Write_Value(wire_16[7:0]), .Output_A(wire_7_1), .Output_B(wire_26_6), .Output());

  wire [0:0] wire_0;
  wire [7:0] wire_1;
  wire [0:0] wire_2;
  wire [7:0] wire_3;
  wire [0:0] wire_4;
  wire [7:0] wire_5;
  wire [7:0] wire_6;
  wire [7:0] wire_7;
  wire [7:0] wire_7_0;
  wire [7:0] wire_7_1;
  wire [7:0] wire_7_2;
  wire [7:0] wire_7_3;
  wire [7:0] wire_7_4;
  wire [7:0] wire_7_5;
  wire [7:0] wire_7_6;
  wire [7:0] wire_7_7;
  assign wire_7 = wire_7_0|wire_7_1|wire_7_2|wire_7_3|wire_7_4|wire_7_5|wire_7_6|wire_7_7;
  wire [7:0] wire_8;
  wire [7:0] wire_8_0;
  wire [7:0] wire_8_1;
  assign wire_8 = wire_8_0|wire_8_1;
  wire [7:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [63:0] wire_16;
  wire [63:0] wire_16_0;
  wire [63:0] wire_16_1;
  wire [63:0] wire_16_2;
  wire [63:0] wire_16_3;
  wire [63:0] wire_16_4;
  wire [63:0] wire_16_5;
  wire [63:0] wire_16_6;
  wire [63:0] wire_16_7;
  wire [63:0] wire_16_8;
  assign wire_16 = wire_16_0|wire_16_1|wire_16_2|wire_16_3|wire_16_4|wire_16_5|wire_16_6|wire_16_7|wire_16_8;
  wire [0:0] wire_17;
  wire [7:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [7:0] wire_26;
  wire [7:0] wire_26_0;
  wire [7:0] wire_26_1;
  wire [7:0] wire_26_2;
  wire [7:0] wire_26_3;
  wire [7:0] wire_26_4;
  wire [7:0] wire_26_5;
  wire [7:0] wire_26_6;
  wire [7:0] wire_26_7;
  assign wire_26 = wire_26_0|wire_26_1|wire_26_2|wire_26_3|wire_26_4|wire_26_5|wire_26_6|wire_26_7;
  wire [0:0] wire_27;
  wire [0:0] wire_27_0;
  wire [0:0] wire_27_1;
  wire [0:0] wire_27_2;
  wire [0:0] wire_27_3;
  wire [0:0] wire_27_4;
  wire [0:0] wire_27_5;
  assign wire_27 = wire_27_0|wire_27_1|wire_27_2|wire_27_3|wire_27_4|wire_27_5;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  assign arch_input_enable = wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [7:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [63:0] wire_42;
  wire [7:0] wire_43;
  wire [0:0] wire_44;
  wire [63:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [7:0] wire_51;
  wire [0:0] wire_52;
  wire [7:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [7:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [7:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;
  wire [7:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  assign arch_output_enable = wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [7:0] wire_80;
  wire [0:0] wire_81;
  wire [63:0] wire_82;
  wire [0:0] wire_83;
  wire [7:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [7:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  wire [7:0] wire_94;
  wire [0:0] wire_95;
  wire [0:0] wire_96;
  wire [0:0] wire_97;
  wire [7:0] wire_98;
  wire [0:0] wire_99;
  wire [0:0] wire_100;
  wire [63:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [0:0] wire_106;
  wire [7:0] wire_107;
  wire [0:0] wire_108;
  wire [0:0] wire_109;
  wire [0:0] wire_110;

endmodule
